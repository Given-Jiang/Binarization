-- Binarization_GN_Binarization_Binarization_Module.vhd

-- Generated using ACDS version 13.1 162 at 2015.02.12.09:18:23

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Binarization_GN_Binarization_Binarization_Module is
	port (
		sop       : in  std_logic                     := '0';             --       sop.wire
		writedata : in  std_logic_vector(31 downto 0) := (others => '0'); -- writedata.wire
		eop       : in  std_logic                     := '0';             --       eop.wire
		addr      : in  std_logic_vector(1 downto 0)  := (others => '0'); --      addr.wire
		write     : in  std_logic                     := '0';             --     write.wire
		Clock     : in  std_logic                     := '0';             --     Clock.clk
		aclr      : in  std_logic                     := '0';             --          .reset
		data_out  : out std_logic_vector(23 downto 0);                    --  data_out.wire
		data_in   : in  std_logic_vector(23 downto 0) := (others => '0')  --   data_in.wire
	);
end entity Binarization_GN_Binarization_Binarization_Module;

architecture rtl of Binarization_GN_Binarization_Binarization_Module is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_cast_GNKXX25S2S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNKXX25S2S;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component alt_dspbuilder_multiplexer_GNCALBUTDR is
		generic (
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0;
			width                  : positive := 8;
			pipeline               : natural  := 0;
			number_inputs          : natural  := 4
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(23 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNCALBUTDR;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_constant_GNZEH3JAKA is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNZEH3JAKA;

	component alt_dspbuilder_port_GN6TDLHAW6 is
		port (
			input  : in  std_logic_vector(1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GN6TDLHAW6;

	component alt_dspbuilder_constant_GNNKZSYI73 is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNNKZSYI73;

	component alt_dspbuilder_constant_GNLMV7GZFA is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNLMV7GZFA;

	component alt_dspbuilder_if_statement_GNYT6HZJI5 is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                       -- wire
			a    : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(7 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GNYT6HZJI5;

	component alt_dspbuilder_delay_GNUECIBFDH is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNUECIBFDH;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V;

	component alt_dspbuilder_decoder_GNSCEXJCJK is
		generic (
			decode   : string  := "00000000";
			pipeline : natural := 0;
			width    : natural := 8
		);
		port (
			aclr  : in  std_logic                          := 'X';             -- clk
			clock : in  std_logic                          := 'X';             -- clk
			data  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			dec   : out std_logic;                                             -- wire
			ena   : in  std_logic                          := 'X';             -- wire
			sclr  : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_decoder_GNSCEXJCJK;

	component alt_dspbuilder_delay_GNVTJPHWYT is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNVTJPHWYT;

	component alt_dspbuilder_if_statement_GN7VA7SRUP is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                        -- wire
			a    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			c    : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GN7VA7SRUP;

	component alt_dspbuilder_delay_GNHYCSAEGT is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNHYCSAEGT;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component alt_dspbuilder_decoder_GNM4LOIHXZ is
		generic (
			decode   : string  := "00000000";
			pipeline : natural := 0;
			width    : natural := 8
		);
		port (
			aclr  : in  std_logic                          := 'X';             -- clk
			clock : in  std_logic                          := 'X';             -- clk
			data  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			dec   : out std_logic;                                             -- wire
			ena   : in  std_logic                          := 'X';             -- wire
			sclr  : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_decoder_GNM4LOIHXZ;

	component alt_dspbuilder_cast_GN7PRGDOVA is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN7PRGDOVA;

	component alt_dspbuilder_cast_GNSB3OXIQS is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			output : out std_logic                                        -- wire
		);
	end component alt_dspbuilder_cast_GNSB3OXIQS;

	component alt_dspbuilder_cast_GN46N4UJ5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic                    := 'X'; -- wire
			output : out std_logic_vector(0 downto 0)         -- wire
		);
	end component alt_dspbuilder_cast_GN46N4UJ5S;

	signal multiplexeruser_aclrgnd_output_wire  : std_logic;                     -- Multiplexeruser_aclrGND:output -> Multiplexer:user_aclr
	signal multiplexerenavcc_output_wire        : std_logic;                     -- MultiplexerenaVCC:output -> Multiplexer:ena
	signal decoder1sclrgnd_output_wire          : std_logic;                     -- Decoder1sclrGND:output -> Decoder1:sclr
	signal decoder1enavcc_output_wire           : std_logic;                     -- Decoder1enaVCC:output -> Decoder1:ena
	signal delay3sclrgnd_output_wire            : std_logic;                     -- Delay3sclrGND:output -> Delay3:sclr
	signal multiplexer1user_aclrgnd_output_wire : std_logic;                     -- Multiplexer1user_aclrGND:output -> Multiplexer1:user_aclr
	signal multiplexer1enavcc_output_wire       : std_logic;                     -- Multiplexer1enaVCC:output -> Multiplexer1:ena
	signal delay1sclrgnd_output_wire            : std_logic;                     -- Delay1sclrGND:output -> Delay1:sclr
	signal delay1enavcc_output_wire             : std_logic;                     -- Delay1enaVCC:output -> Delay1:ena
	signal delay2sclrgnd_output_wire            : std_logic;                     -- Delay2sclrGND:output -> Delay2:sclr
	signal decodersclrgnd_output_wire           : std_logic;                     -- DecodersclrGND:output -> Decoder:sclr
	signal decoderenavcc_output_wire            : std_logic;                     -- DecoderenaVCC:output -> Decoder:ena
	signal addr_0_output_wire                   : std_logic_vector(1 downto 0);  -- addr_0:output -> Decoder:data
	signal bus_conversion1_output_wire          : std_logic_vector(7 downto 0);  -- Bus_Conversion1:output -> Delay2:input
	signal delay2_output_wire                   : std_logic_vector(7 downto 0);  -- Delay2:output -> Delay3:input
	signal data_in_0_output_wire                : std_logic_vector(23 downto 0); -- data_in_0:output -> [Bus_Conversion:input, Decoder1:data, If_Statement1:a, Multiplexer:in0]
	signal bus_conversion_output_wire           : std_logic_vector(7 downto 0);  -- Bus_Conversion:output -> If_Statement:a
	signal delay3_output_wire                   : std_logic_vector(7 downto 0);  -- Delay3:output -> If_Statement:b
	signal constant3_output_wire                : std_logic_vector(23 downto 0); -- Constant3:output -> If_Statement1:b
	signal constant4_output_wire                : std_logic_vector(23 downto 0); -- Constant4:output -> If_Statement1:c
	signal if_statement1_true_wire              : std_logic;                     -- If_Statement1:true -> Logical_Bit_Operator:data0
	signal sop_0_output_wire                    : std_logic;                     -- sop_0:output -> [Logical_Bit_Operator3:data0, Logical_Bit_Operator:data1]
	signal logical_bit_operator_result_wire     : std_logic;                     -- Logical_Bit_Operator:result -> [Delay:ena, cast2:input]
	signal eop_0_output_wire                    : std_logic;                     -- eop_0:output -> Logical_Bit_Operator1:data0
	signal decoder_dec_wire                     : std_logic;                     -- Decoder:dec -> Logical_Bit_Operator2:data0
	signal write_0_output_wire                  : std_logic;                     -- write_0:output -> Logical_Bit_Operator2:data1
	signal logical_bit_operator2_result_wire    : std_logic;                     -- Logical_Bit_Operator2:result -> Delay2:ena
	signal decoder1_dec_wire                    : std_logic;                     -- Decoder1:dec -> Logical_Bit_Operator3:data1
	signal logical_bit_operator3_result_wire    : std_logic;                     -- Logical_Bit_Operator3:result -> Delay3:ena
	signal delay_output_wire                    : std_logic_vector(0 downto 0);  -- Delay:output -> [Multiplexer:sel, cast3:input]
	signal constant1_output_wire                : std_logic_vector(23 downto 0); -- Constant1:output -> Multiplexer1:in0
	signal constant2_output_wire                : std_logic_vector(23 downto 0); -- Constant2:output -> Multiplexer1:in1
	signal multiplexer1_result_wire             : std_logic_vector(23 downto 0); -- Multiplexer1:result -> Multiplexer:in1
	signal multiplexer_result_wire              : std_logic_vector(23 downto 0); -- Multiplexer:result -> data_out_0:input
	signal writedata_0_output_wire              : std_logic_vector(31 downto 0); -- writedata_0:output -> cast0:input
	signal cast0_output_wire                    : std_logic_vector(23 downto 0); -- cast0:output -> Bus_Conversion1:input
	signal delay1_output_wire                   : std_logic_vector(0 downto 0);  -- Delay1:output -> cast1:input
	signal cast1_output_wire                    : std_logic;                     -- cast1:output -> Delay:sclr
	signal cast2_output_wire                    : std_logic_vector(0 downto 0);  -- cast2:output -> Delay:input
	signal cast3_output_wire                    : std_logic;                     -- cast3:output -> Logical_Bit_Operator1:data1
	signal logical_bit_operator1_result_wire    : std_logic;                     -- Logical_Bit_Operator1:result -> cast4:input
	signal cast4_output_wire                    : std_logic_vector(0 downto 0);  -- cast4:output -> Delay1:input
	signal if_statement_true_wire               : std_logic;                     -- If_Statement:true -> cast5:input
	signal cast5_output_wire                    : std_logic_vector(0 downto 0);  -- cast5:output -> Multiplexer1:sel
	signal clock_0_clock_output_reset           : std_logic;                     -- Clock_0:aclr_out -> [Decoder1:aclr, Decoder:aclr, Delay1:aclr, Delay2:aclr, Delay3:aclr, Delay:aclr, Multiplexer1:aclr, Multiplexer:aclr]
	signal clock_0_clock_output_clk             : std_logic;                     -- Clock_0:clock_out -> [Decoder1:clock, Decoder:clock, Delay1:clock, Delay2:clock, Delay3:clock, Delay:clock, Multiplexer1:clock, Multiplexer:clock]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	bus_conversion1 : component alt_dspbuilder_cast_GNKXX25S2S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast0_output_wire,           --  input.wire
			output => bus_conversion1_output_wire  -- output.wire
		);

	writedata_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => writedata,               --  input.wire
			output => writedata_0_output_wire  -- output.wire
		);

	multiplexer : component alt_dspbuilder_multiplexer_GNCALBUTDR
		generic map (
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0,
			width                  => 24,
			pipeline               => 0,
			number_inputs          => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			sel       => delay_output_wire,                   --        sel.wire
			result    => multiplexer_result_wire,             --     result.wire
			ena       => multiplexerenavcc_output_wire,       --        ena.wire
			user_aclr => multiplexeruser_aclrgnd_output_wire, --  user_aclr.wire
			in0       => data_in_0_output_wire,               --        in0.wire
			in1       => multiplexer1_result_wire             --        in1.wire
		);

	multiplexeruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexeruser_aclrgnd_output_wire  -- output.wire
		);

	multiplexerenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexerenavcc_output_wire  -- output.wire
		);

	bus_conversion : component alt_dspbuilder_cast_GNKXX25S2S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_in_0_output_wire,      --  input.wire
			output => bus_conversion_output_wire  -- output.wire
		);

	constant4 : component alt_dspbuilder_constant_GNZEH3JAKA
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000001111",
			width      => 24
		)
		port map (
			output => constant4_output_wire  -- output.wire
		);

	addr_0 : component alt_dspbuilder_port_GN6TDLHAW6
		port map (
			input  => addr,               --  input.wire
			output => addr_0_output_wire  -- output.wire
		);

	constant3 : component alt_dspbuilder_constant_GNNKZSYI73
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000000000",
			width      => 24
		)
		port map (
			output => constant3_output_wire  -- output.wire
		);

	constant2 : component alt_dspbuilder_constant_GNLMV7GZFA
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "111111111111111111111111",
			width      => 24
		)
		port map (
			output => constant2_output_wire  -- output.wire
		);

	if_statement : component alt_dspbuilder_if_statement_GNYT6HZJI5
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "a>b",
			number_inputs   => 2,
			width           => 8
		)
		port map (
			true => if_statement_true_wire,     -- true.wire
			a    => bus_conversion_output_wire, --    a.wire
			b    => delay3_output_wire          --    b.wire
		);

	constant1 : component alt_dspbuilder_constant_GNNKZSYI73
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000000000",
			width      => 24
		)
		port map (
			output => constant1_output_wire  -- output.wire
		);

	delay : component alt_dspbuilder_delay_GNUECIBFDH
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "0",
			width      => 1
		)
		port map (
			input  => cast2_output_wire,                --      input.wire
			clock  => clock_0_clock_output_clk,         -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,       --           .reset
			output => delay_output_wire,                --     output.wire
			sclr   => cast1_output_wire,                --       sclr.wire
			ena    => logical_bit_operator_result_wire  --        ena.wire
		);

	write_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => write,               --  input.wire
			output => write_0_output_wire  -- output.wire
		);

	logical_bit_operator3 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator3_result_wire, -- result.wire
			data0  => sop_0_output_wire,                 --  data0.wire
			data1  => decoder1_dec_wire                  --  data1.wire
		);

	eop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => eop,               --  input.wire
			output => eop_0_output_wire  -- output.wire
		);

	logical_bit_operator2 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator2_result_wire, -- result.wire
			data0  => decoder_dec_wire,                  --  data0.wire
			data1  => write_0_output_wire                --  data1.wire
		);

	logical_bit_operator1 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator1_result_wire, -- result.wire
			data0  => eop_0_output_wire,                 --  data0.wire
			data1  => cast3_output_wire                  --  data1.wire
		);

	decoder1 : component alt_dspbuilder_decoder_GNSCEXJCJK
		generic map (
			decode   => "000000000000000000001111",
			pipeline => 0,
			width    => 24
		)
		port map (
			clock => clock_0_clock_output_clk,    -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,  --           .reset
			data  => data_in_0_output_wire,       --       data.wire
			dec   => decoder1_dec_wire,           --        dec.wire
			sclr  => decoder1sclrgnd_output_wire, --       sclr.wire
			ena   => decoder1enavcc_output_wire   --        ena.wire
		);

	decoder1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decoder1sclrgnd_output_wire  -- output.wire
		);

	decoder1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoder1enavcc_output_wire  -- output.wire
		);

	logical_bit_operator : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator_result_wire, -- result.wire
			data0  => if_statement1_true_wire,          --  data0.wire
			data1  => sop_0_output_wire                 --  data1.wire
		);

	delay3 : component alt_dspbuilder_delay_GNVTJPHWYT
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "01111111",
			width      => 8
		)
		port map (
			input  => delay2_output_wire,                --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay3_output_wire,                --     output.wire
			sclr   => delay3sclrgnd_output_wire,         --       sclr.wire
			ena    => logical_bit_operator3_result_wire  --        ena.wire
		);

	delay3sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay3sclrgnd_output_wire  -- output.wire
		);

	if_statement1 : component alt_dspbuilder_if_statement_GN7VA7SRUP
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "(a=b) and (a /= c)",
			number_inputs   => 3,
			width           => 24
		)
		port map (
			true => if_statement1_true_wire, -- true.wire
			a    => data_in_0_output_wire,   --    a.wire
			b    => constant3_output_wire,   --    b.wire
			c    => constant4_output_wire    --    c.wire
		);

	sop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sop,               --  input.wire
			output => sop_0_output_wire  -- output.wire
		);

	multiplexer1 : component alt_dspbuilder_multiplexer_GNCALBUTDR
		generic map (
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0,
			width                  => 24,
			pipeline               => 0,
			number_inputs          => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast5_output_wire,                    --        sel.wire
			result    => multiplexer1_result_wire,             --     result.wire
			ena       => multiplexer1enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer1user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => constant1_output_wire,                --        in0.wire
			in1       => constant2_output_wire                 --        in1.wire
		);

	multiplexer1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer1user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer1enavcc_output_wire  -- output.wire
		);

	delay1 : component alt_dspbuilder_delay_GNHYCSAEGT
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 0,
			BitPattern => "0",
			width      => 1
		)
		port map (
			input  => cast4_output_wire,          --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay1_output_wire,         --     output.wire
			sclr   => delay1sclrgnd_output_wire,  --       sclr.wire
			ena    => delay1enavcc_output_wire    --        ena.wire
		);

	delay1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay1sclrgnd_output_wire  -- output.wire
		);

	delay1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delay1enavcc_output_wire  -- output.wire
		);

	delay2 : component alt_dspbuilder_delay_GNVTJPHWYT
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "01111111",
			width      => 8
		)
		port map (
			input  => bus_conversion1_output_wire,       --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay2_output_wire,                --     output.wire
			sclr   => delay2sclrgnd_output_wire,         --       sclr.wire
			ena    => logical_bit_operator2_result_wire  --        ena.wire
		);

	delay2sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay2sclrgnd_output_wire  -- output.wire
		);

	data_out_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => multiplexer_result_wire, --  input.wire
			output => data_out                 -- output.wire
		);

	data_in_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => data_in,               --  input.wire
			output => data_in_0_output_wire  -- output.wire
		);

	decoder : component alt_dspbuilder_decoder_GNM4LOIHXZ
		generic map (
			decode   => "01",
			pipeline => 1,
			width    => 2
		)
		port map (
			clock => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset, --           .reset
			data  => addr_0_output_wire,         --       data.wire
			dec   => decoder_dec_wire,           --        dec.wire
			sclr  => decodersclrgnd_output_wire, --       sclr.wire
			ena   => decoderenavcc_output_wire   --        ena.wire
		);

	decodersclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decodersclrgnd_output_wire  -- output.wire
		);

	decoderenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoderenavcc_output_wire  -- output.wire
		);

	cast0 : component alt_dspbuilder_cast_GN7PRGDOVA
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => writedata_0_output_wire, --  input.wire
			output => cast0_output_wire        -- output.wire
		);

	cast1 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire, --  input.wire
			output => cast1_output_wire   -- output.wire
		);

	cast2 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => logical_bit_operator_result_wire, --  input.wire
			output => cast2_output_wire                 -- output.wire
		);

	cast3 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay_output_wire, --  input.wire
			output => cast3_output_wire  -- output.wire
		);

	cast4 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => logical_bit_operator1_result_wire, --  input.wire
			output => cast4_output_wire                  -- output.wire
		);

	cast5 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => if_statement_true_wire, --  input.wire
			output => cast5_output_wire       -- output.wire
		);

end architecture rtl; -- of Binarization_GN_Binarization_Binarization_Module
